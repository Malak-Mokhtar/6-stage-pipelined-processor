LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY Reg_file IS
    PORT (
        clock
    );
END Reg_file;

ARCHITECTURE arch OF Reg_file IS

BEGIN

END ARCHITECTURE;